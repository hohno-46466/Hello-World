/*
  Verilog HDL
*/

module main();
    initial $display("Hello, World!");
endmodule

// This line also can be a comment line
